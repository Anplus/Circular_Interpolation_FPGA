
module sel_in(	// system connections
				sys_rst_l,
				sys_clk,

				// sync input
				change_readyH

				// data input
				shape,		//1bit
				method,		//2bits
				
				);

always @(change) begin

end


endmodule
