module speed_cal(
);

endmodule
