
module select_out(

		);

endmodule
