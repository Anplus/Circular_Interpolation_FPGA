library verilog;
use verilog.vl_types.all;
entity work_test is
end work_test;
